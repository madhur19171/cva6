module ariane_testharness_wrapper(
    input  logic                           clk_i,
    input  logic                           rtc_i,
    input  logic                           rst_ni,
    output logic [31:0]                    exit_o
);

    wire [63 : 0]   Router_data_out     [1 : 0];
    wire            Router_valid_out    [1 : 0];
    wire            Router_ready_out    [1 : 0];

    wire [63 : 0]   Router_data_in      [1 : 0];
    wire            Router_valid_in     [1 : 0];
    wire            Router_ready_in     [1 : 0];

    ariane_testharness #(.hart_id_in(0)) i_ariane_testharness_0
        (
            .clk_i(clk_i),
            .rtc_i(rtc_i),
            .rst_ni(rst_ni),
            .exit_o(),

            .data_in(Router_data_out[0]), .valid_in(Router_valid_out[0]), .ready_in(Router_ready_out[0]),
            .data_out(Router_data_in[0]), .valid_out(Router_valid_in[0]), .ready_out(Router_ready_in[0])

        );

    ariane_testharness #(.hart_id_in(0)) i_ariane_testharness_1
        (
            .clk_i(clk_i),
            .rtc_i(rtc_i),
            .rst_ni(rst_ni),
            .exit_o(),

            .data_in(Router_data_out[1]), .valid_in(Router_valid_out[1]), .ready_in(Router_ready_out[1]),
            .data_out(Router_data_in[1]), .valid_out(Router_valid_in[1]), .ready_out(Router_ready_in[1])

        );

    Mesh22 mesh22 (
    .clk(clk_i), .rst(~rst_ni),
    .Node0_data_in(Router_data_in[0]), .Node0_valid_in(Router_valid_in[0]), .Node0_ready_in(Router_ready_in[0]),
    .Node0_data_out(Router_data_out[0]), .Node0_valid_out(Router_valid_out[0]), .Node0_ready_out(Router_ready_out[0]),

    .Node1_data_in(), .Node1_valid_in(), .Node1_ready_in(),
    .Node1_data_out(), .Node1_valid_out(), .Node1_ready_out(1),

    .Node2_data_in(), .Node2_valid_in(), .Node2_ready_in(),
    .Node2_data_out(), .Node2_valid_out(), .Node2_ready_out(1),

    .Node3_data_in(Router_data_in[1]), .Node3_valid_in(Router_valid_in[1]), .Node3_ready_in(Router_ready_in[1]),
    .Node3_data_out(Router_data_out[1]), .Node3_valid_out(Router_valid_out[1]), .Node3_ready_out(Router_ready_out[1])
  );
    
endmodule